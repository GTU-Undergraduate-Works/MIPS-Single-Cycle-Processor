module ALU_testbench();



reg [31:0] data1, data2;
reg [3:0] ALUOp;
reg [4:0] shamt;
wire [31:0] result;
wire zero;

ALU opeartionresult(data1, data2, ALUOp, shamt, result, zero);



initial begin

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // ADD
ALUOp = 4'b0001; shamt = 5'b00000; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // AND
ALUOp = 4'b0010; shamt = 5'b00000; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // NOR
ALUOp = 4'b0011; shamt = 5'b00000; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // OR
ALUOp = 4'b0100; shamt = 5'b00000; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // SLL
ALUOp = 4'b0101; shamt = 5'b00010; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // SRL
ALUOp = 4'b0110; shamt = 5'b00011; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // SLT
ALUOp = 4'b0111; shamt = 5'b00011; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // SLTU
ALUOp = 4'b1000; shamt = 5'b00011; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // SUB
ALUOp = 4'b1001; shamt = 5'b00011; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b00000000000000111111111111110000; // SUBU
ALUOp = 4'b1010; shamt = 5'b00011; #20;

data1 = 32'b10000001010101010101111111001101; data2 = 32'b10000001010101010101111111001101; // SUB
ALUOp = 4'b1001; shamt = 5'b00011; #20;

data1 = 32'b00000000000000111111111111110000; data2 = 32'b00000000000000111111111111110000; // SUBU
ALUOp = 4'b1010; shamt = 5'b00011; #20;

end

initial begin
	$monitor("time = %2d\nALUOp = %4b\nshamt = %5b\ndata1 =  %32b\ndata2 =  %32b\nresult = %32b\nzero = %1b\n\n",
				$time, ALUOp, shamt, data1, data2, result, zero);
end


endmodule
